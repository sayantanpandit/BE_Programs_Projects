----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:13:36 03/29/2016 
-- Design Name: 
-- Module Name:    JK_FF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity JK_FF is
    Port ( J : in  STD_LOGIC;
           K : in  STD_LOGIC;
           CLOCK : in  STD_LOGIC;
           Q : out  STD_LOGIC;
           QB : out  STD_LOGIC);
end JK_FF;

architecture Behavioral of JK_FF is
begin
	PROCESS(CLOCK)
	variable TMP: std_logic;
	begin
		if(CLOCK='1' and CLOCK'EVENT) then
						if(J='0' and K='0')then
								TMP:=TMP;
						elsif(J='1' and K='1')then
								TMP:= not TMP;
						elsif(J='0' and K='1')then
								TMP:='0';
						else
								TMP:='1';
						end if;
		end if;
		Q<=TMP;
		QB<=not TMP;
end PROCESS;
end Behavioral;

