module segment(D,C,B,A,a,b,c,d,e,f,g);

input D,C,B,A;
output a,b,c,d,e,f,g;

assign a = ((!D)&(!C)&(!B)&(!A)) | ((!D)&(!C)&(B)&(!A)) | ((!D)&(!C)&(B)&(A)) | ((!D)&(C)&(!B)&(A)) | ((!D)&(C)&(B)&(A)) | ((D)&(!C)&(!B)&(!A)) | ((D)&(!C)&(!B)&(A));
assign b = ((!D)&(!C)&(!B)&(!A)) | ((!D)&(!C)&(!B)&(A)) | ((!D)&(!C)&(B)&(!A)) | ((!D)&(!C)&(B)&(A)) | ((!D)&(C)&(!B)&(!A)) | ((!D)&(C)&(B)&(A)) | ((D)&(!C)&(!B)&(!A)) | ((D)&(!C)&(!B)&(A));
assign c = ((!D)&(!C)&(!B)&(!A)) | ((!D)&(!C)&(!B)&(A)) | ((!D)&(!C)&(B)&(A)) | ((!D)&(C)&(!B)&(!A)) | ((!D)&(C)&(!B)&(A)) | ((!D)&(C)&(B)&(!A)) | ((!D)&(C)&(B)&(A)) | ((D)&(!C)&(!B)&(!A)) | ((D)&(!C)&(!B)&(A));
assign d = ((!D)&(!C)&(!B)&(!A)) | ((!D)&(!C)&(B)&(!A)) | ((!D)&(!C)&(B)&(A)) | ((!D)&(C)&(!B)&(A)) | ((!D)&(C)&(B)&(!A)) | ((D)&(!C)&(!B)&(!A));
assign e = ((!D)&(!C)&(!B)&(!A)) | ((!D)&(!C)&(B)&(!A)) | ((!D)&(C)&(B)&(!A)) | ((D)&(!C)&(!B)&(!A));
assign f = ((!D)&(!C)&(!B)&(!A)) | ((!D)&(C)&(!B)&(!A)) | ((!D)&(C)&(!B)&(A)) | ((!D)&(C)&(B)&(!A)) | ((D)&(!C)&(!B)&(!A)) | ((D)&(!C)&(!B)&(A));
assign g = ((!D)&(!C)&(B)&(!A)) | ((!D)&(!C)&(B)&(A)) | ((!D)&(C)&(!B)&(!A)) | ((!D)&(C)&(!B)&(A)) | ((!D)&(C)&(B)&(!A)) | ((D)&(!C)&(!B)&(!A)) | ((D)&(!C)&(!B)&(A));

endmodule